library ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
ENTITY Preprocessor IS
	PORT(clk: IN STD_LOGIC;
		  reset : IN STD_LOGIC;
		  ready : IN STD_LOGIC;
		  readyBlock:IN STD_LOGIC;
		  lastBlock:OUT STD_LOGIC;
		  --xzeros:out std_logic_vector(0 to 63);
		  k,n: out integer;
		  --a1:out unsigned(0 to 63);
		  --a2:out unsigned(0 to 63);
		  --messageString : IN string:="ab";
		  --lengthInteger:out integer;
		  --out1:OUT std_logic_vector(0 to 15);
		  messageBit : OUT std_logic_vector(0 to 511)
		  --messsageLenVecotr : out std_LOGIC_VECTOR(0 to 63)
		 );
end Preprocessor;

ARCHITECTURE behavioral of Preprocessor IS
	--signal input : string(1 to 2);
	constant ss : string :="abcdefghijklmnopqrstuvwxyzabcdefghijklmnopqrstuvwxyzabcd";
	signal output:std_logic_vector(0 to ss'length*8 +(447- ss'length*8) mod 512+64);
	signal messageLength : std_LOGIC_VECTOR(0 to 63);
	signal len_unsigned,k0 : unsigned (0 to 63);
	signal nBlocks,x:integer;
	
	
	begin
		PROCESS(clk,ready,readyBlock)
		begin	
			if(clk'Event and clk='1' and ready ='1')then
				k<=output'length;
				nBlocks<=output'length/512;
				IF(nBlocks /= 0)then
					x<=1;
				end if;
				n<=nBlocks;
				len_unsigned<=shift_left(to_unsigned(ss'length,64),3);
				messageLength<= std_logic_vector(len_unsigned);

				k0<=(447- len_unsigned) mod 512;			
				
				output(TO_INTEGER(len_unsigned))<='1';
				
				for i in 1 to 447 loop
					exit when i=((TO_INTEGER(k0))+1);
					output((TO_INTEGER(len_unsigned)) +i)<='0'; 
				end loop;
				
				
				for i in  ss'range loop
					output((8*i)-8 to (8*i)-1)<=std_logic_vector(to_unsigned(character'pos(ss(i)),8));
				end loop;
								
				output(448 to 511)<=messageLength;

			elsif(clk'Event and clk='1' and ready='0')then
				output<=std_logic_vector(to_unsigned(0,output'length));
			elsif(clk'Event and clk='1' and readyBlock='0')then
				if(x=nBlocks)then
					lastBlock<='1';
					x<=0;
				else
					x<=x+1;
				end if;
			end if;
		end process;
			messageBit<=output(x*512 to x*512+511);
end behavioral;