library verilog;
use verilog.vl_types.all;
entity MessageScheduler is
    port(
        clk             : in     vl_logic;
        M               : in     vl_logic_vector(511 downto 0);
        W_63_0          : out    vl_logic;
        W_63_1          : out    vl_logic;
        W_63_2          : out    vl_logic;
        W_63_3          : out    vl_logic;
        W_63_4          : out    vl_logic;
        W_63_5          : out    vl_logic;
        W_63_6          : out    vl_logic;
        W_63_7          : out    vl_logic;
        W_63_8          : out    vl_logic;
        W_63_9          : out    vl_logic;
        W_63_10         : out    vl_logic;
        W_63_11         : out    vl_logic;
        W_63_12         : out    vl_logic;
        W_63_13         : out    vl_logic;
        W_63_14         : out    vl_logic;
        W_63_15         : out    vl_logic;
        W_63_16         : out    vl_logic;
        W_63_17         : out    vl_logic;
        W_63_18         : out    vl_logic;
        W_63_19         : out    vl_logic;
        W_63_20         : out    vl_logic;
        W_63_21         : out    vl_logic;
        W_63_22         : out    vl_logic;
        W_63_23         : out    vl_logic;
        W_63_24         : out    vl_logic;
        W_63_25         : out    vl_logic;
        W_63_26         : out    vl_logic;
        W_63_27         : out    vl_logic;
        W_63_28         : out    vl_logic;
        W_63_29         : out    vl_logic;
        W_63_30         : out    vl_logic;
        W_63_31         : out    vl_logic;
        W_62_0          : out    vl_logic;
        W_62_1          : out    vl_logic;
        W_62_2          : out    vl_logic;
        W_62_3          : out    vl_logic;
        W_62_4          : out    vl_logic;
        W_62_5          : out    vl_logic;
        W_62_6          : out    vl_logic;
        W_62_7          : out    vl_logic;
        W_62_8          : out    vl_logic;
        W_62_9          : out    vl_logic;
        W_62_10         : out    vl_logic;
        W_62_11         : out    vl_logic;
        W_62_12         : out    vl_logic;
        W_62_13         : out    vl_logic;
        W_62_14         : out    vl_logic;
        W_62_15         : out    vl_logic;
        W_62_16         : out    vl_logic;
        W_62_17         : out    vl_logic;
        W_62_18         : out    vl_logic;
        W_62_19         : out    vl_logic;
        W_62_20         : out    vl_logic;
        W_62_21         : out    vl_logic;
        W_62_22         : out    vl_logic;
        W_62_23         : out    vl_logic;
        W_62_24         : out    vl_logic;
        W_62_25         : out    vl_logic;
        W_62_26         : out    vl_logic;
        W_62_27         : out    vl_logic;
        W_62_28         : out    vl_logic;
        W_62_29         : out    vl_logic;
        W_62_30         : out    vl_logic;
        W_62_31         : out    vl_logic;
        W_61_0          : out    vl_logic;
        W_61_1          : out    vl_logic;
        W_61_2          : out    vl_logic;
        W_61_3          : out    vl_logic;
        W_61_4          : out    vl_logic;
        W_61_5          : out    vl_logic;
        W_61_6          : out    vl_logic;
        W_61_7          : out    vl_logic;
        W_61_8          : out    vl_logic;
        W_61_9          : out    vl_logic;
        W_61_10         : out    vl_logic;
        W_61_11         : out    vl_logic;
        W_61_12         : out    vl_logic;
        W_61_13         : out    vl_logic;
        W_61_14         : out    vl_logic;
        W_61_15         : out    vl_logic;
        W_61_16         : out    vl_logic;
        W_61_17         : out    vl_logic;
        W_61_18         : out    vl_logic;
        W_61_19         : out    vl_logic;
        W_61_20         : out    vl_logic;
        W_61_21         : out    vl_logic;
        W_61_22         : out    vl_logic;
        W_61_23         : out    vl_logic;
        W_61_24         : out    vl_logic;
        W_61_25         : out    vl_logic;
        W_61_26         : out    vl_logic;
        W_61_27         : out    vl_logic;
        W_61_28         : out    vl_logic;
        W_61_29         : out    vl_logic;
        W_61_30         : out    vl_logic;
        W_61_31         : out    vl_logic;
        W_60_0          : out    vl_logic;
        W_60_1          : out    vl_logic;
        W_60_2          : out    vl_logic;
        W_60_3          : out    vl_logic;
        W_60_4          : out    vl_logic;
        W_60_5          : out    vl_logic;
        W_60_6          : out    vl_logic;
        W_60_7          : out    vl_logic;
        W_60_8          : out    vl_logic;
        W_60_9          : out    vl_logic;
        W_60_10         : out    vl_logic;
        W_60_11         : out    vl_logic;
        W_60_12         : out    vl_logic;
        W_60_13         : out    vl_logic;
        W_60_14         : out    vl_logic;
        W_60_15         : out    vl_logic;
        W_60_16         : out    vl_logic;
        W_60_17         : out    vl_logic;
        W_60_18         : out    vl_logic;
        W_60_19         : out    vl_logic;
        W_60_20         : out    vl_logic;
        W_60_21         : out    vl_logic;
        W_60_22         : out    vl_logic;
        W_60_23         : out    vl_logic;
        W_60_24         : out    vl_logic;
        W_60_25         : out    vl_logic;
        W_60_26         : out    vl_logic;
        W_60_27         : out    vl_logic;
        W_60_28         : out    vl_logic;
        W_60_29         : out    vl_logic;
        W_60_30         : out    vl_logic;
        W_60_31         : out    vl_logic;
        W_59_0          : out    vl_logic;
        W_59_1          : out    vl_logic;
        W_59_2          : out    vl_logic;
        W_59_3          : out    vl_logic;
        W_59_4          : out    vl_logic;
        W_59_5          : out    vl_logic;
        W_59_6          : out    vl_logic;
        W_59_7          : out    vl_logic;
        W_59_8          : out    vl_logic;
        W_59_9          : out    vl_logic;
        W_59_10         : out    vl_logic;
        W_59_11         : out    vl_logic;
        W_59_12         : out    vl_logic;
        W_59_13         : out    vl_logic;
        W_59_14         : out    vl_logic;
        W_59_15         : out    vl_logic;
        W_59_16         : out    vl_logic;
        W_59_17         : out    vl_logic;
        W_59_18         : out    vl_logic;
        W_59_19         : out    vl_logic;
        W_59_20         : out    vl_logic;
        W_59_21         : out    vl_logic;
        W_59_22         : out    vl_logic;
        W_59_23         : out    vl_logic;
        W_59_24         : out    vl_logic;
        W_59_25         : out    vl_logic;
        W_59_26         : out    vl_logic;
        W_59_27         : out    vl_logic;
        W_59_28         : out    vl_logic;
        W_59_29         : out    vl_logic;
        W_59_30         : out    vl_logic;
        W_59_31         : out    vl_logic;
        W_58_0          : out    vl_logic;
        W_58_1          : out    vl_logic;
        W_58_2          : out    vl_logic;
        W_58_3          : out    vl_logic;
        W_58_4          : out    vl_logic;
        W_58_5          : out    vl_logic;
        W_58_6          : out    vl_logic;
        W_58_7          : out    vl_logic;
        W_58_8          : out    vl_logic;
        W_58_9          : out    vl_logic;
        W_58_10         : out    vl_logic;
        W_58_11         : out    vl_logic;
        W_58_12         : out    vl_logic;
        W_58_13         : out    vl_logic;
        W_58_14         : out    vl_logic;
        W_58_15         : out    vl_logic;
        W_58_16         : out    vl_logic;
        W_58_17         : out    vl_logic;
        W_58_18         : out    vl_logic;
        W_58_19         : out    vl_logic;
        W_58_20         : out    vl_logic;
        W_58_21         : out    vl_logic;
        W_58_22         : out    vl_logic;
        W_58_23         : out    vl_logic;
        W_58_24         : out    vl_logic;
        W_58_25         : out    vl_logic;
        W_58_26         : out    vl_logic;
        W_58_27         : out    vl_logic;
        W_58_28         : out    vl_logic;
        W_58_29         : out    vl_logic;
        W_58_30         : out    vl_logic;
        W_58_31         : out    vl_logic;
        W_57_0          : out    vl_logic;
        W_57_1          : out    vl_logic;
        W_57_2          : out    vl_logic;
        W_57_3          : out    vl_logic;
        W_57_4          : out    vl_logic;
        W_57_5          : out    vl_logic;
        W_57_6          : out    vl_logic;
        W_57_7          : out    vl_logic;
        W_57_8          : out    vl_logic;
        W_57_9          : out    vl_logic;
        W_57_10         : out    vl_logic;
        W_57_11         : out    vl_logic;
        W_57_12         : out    vl_logic;
        W_57_13         : out    vl_logic;
        W_57_14         : out    vl_logic;
        W_57_15         : out    vl_logic;
        W_57_16         : out    vl_logic;
        W_57_17         : out    vl_logic;
        W_57_18         : out    vl_logic;
        W_57_19         : out    vl_logic;
        W_57_20         : out    vl_logic;
        W_57_21         : out    vl_logic;
        W_57_22         : out    vl_logic;
        W_57_23         : out    vl_logic;
        W_57_24         : out    vl_logic;
        W_57_25         : out    vl_logic;
        W_57_26         : out    vl_logic;
        W_57_27         : out    vl_logic;
        W_57_28         : out    vl_logic;
        W_57_29         : out    vl_logic;
        W_57_30         : out    vl_logic;
        W_57_31         : out    vl_logic;
        W_56_0          : out    vl_logic;
        W_56_1          : out    vl_logic;
        W_56_2          : out    vl_logic;
        W_56_3          : out    vl_logic;
        W_56_4          : out    vl_logic;
        W_56_5          : out    vl_logic;
        W_56_6          : out    vl_logic;
        W_56_7          : out    vl_logic;
        W_56_8          : out    vl_logic;
        W_56_9          : out    vl_logic;
        W_56_10         : out    vl_logic;
        W_56_11         : out    vl_logic;
        W_56_12         : out    vl_logic;
        W_56_13         : out    vl_logic;
        W_56_14         : out    vl_logic;
        W_56_15         : out    vl_logic;
        W_56_16         : out    vl_logic;
        W_56_17         : out    vl_logic;
        W_56_18         : out    vl_logic;
        W_56_19         : out    vl_logic;
        W_56_20         : out    vl_logic;
        W_56_21         : out    vl_logic;
        W_56_22         : out    vl_logic;
        W_56_23         : out    vl_logic;
        W_56_24         : out    vl_logic;
        W_56_25         : out    vl_logic;
        W_56_26         : out    vl_logic;
        W_56_27         : out    vl_logic;
        W_56_28         : out    vl_logic;
        W_56_29         : out    vl_logic;
        W_56_30         : out    vl_logic;
        W_56_31         : out    vl_logic;
        W_55_0          : out    vl_logic;
        W_55_1          : out    vl_logic;
        W_55_2          : out    vl_logic;
        W_55_3          : out    vl_logic;
        W_55_4          : out    vl_logic;
        W_55_5          : out    vl_logic;
        W_55_6          : out    vl_logic;
        W_55_7          : out    vl_logic;
        W_55_8          : out    vl_logic;
        W_55_9          : out    vl_logic;
        W_55_10         : out    vl_logic;
        W_55_11         : out    vl_logic;
        W_55_12         : out    vl_logic;
        W_55_13         : out    vl_logic;
        W_55_14         : out    vl_logic;
        W_55_15         : out    vl_logic;
        W_55_16         : out    vl_logic;
        W_55_17         : out    vl_logic;
        W_55_18         : out    vl_logic;
        W_55_19         : out    vl_logic;
        W_55_20         : out    vl_logic;
        W_55_21         : out    vl_logic;
        W_55_22         : out    vl_logic;
        W_55_23         : out    vl_logic;
        W_55_24         : out    vl_logic;
        W_55_25         : out    vl_logic;
        W_55_26         : out    vl_logic;
        W_55_27         : out    vl_logic;
        W_55_28         : out    vl_logic;
        W_55_29         : out    vl_logic;
        W_55_30         : out    vl_logic;
        W_55_31         : out    vl_logic;
        W_54_0          : out    vl_logic;
        W_54_1          : out    vl_logic;
        W_54_2          : out    vl_logic;
        W_54_3          : out    vl_logic;
        W_54_4          : out    vl_logic;
        W_54_5          : out    vl_logic;
        W_54_6          : out    vl_logic;
        W_54_7          : out    vl_logic;
        W_54_8          : out    vl_logic;
        W_54_9          : out    vl_logic;
        W_54_10         : out    vl_logic;
        W_54_11         : out    vl_logic;
        W_54_12         : out    vl_logic;
        W_54_13         : out    vl_logic;
        W_54_14         : out    vl_logic;
        W_54_15         : out    vl_logic;
        W_54_16         : out    vl_logic;
        W_54_17         : out    vl_logic;
        W_54_18         : out    vl_logic;
        W_54_19         : out    vl_logic;
        W_54_20         : out    vl_logic;
        W_54_21         : out    vl_logic;
        W_54_22         : out    vl_logic;
        W_54_23         : out    vl_logic;
        W_54_24         : out    vl_logic;
        W_54_25         : out    vl_logic;
        W_54_26         : out    vl_logic;
        W_54_27         : out    vl_logic;
        W_54_28         : out    vl_logic;
        W_54_29         : out    vl_logic;
        W_54_30         : out    vl_logic;
        W_54_31         : out    vl_logic;
        W_53_0          : out    vl_logic;
        W_53_1          : out    vl_logic;
        W_53_2          : out    vl_logic;
        W_53_3          : out    vl_logic;
        W_53_4          : out    vl_logic;
        W_53_5          : out    vl_logic;
        W_53_6          : out    vl_logic;
        W_53_7          : out    vl_logic;
        W_53_8          : out    vl_logic;
        W_53_9          : out    vl_logic;
        W_53_10         : out    vl_logic;
        W_53_11         : out    vl_logic;
        W_53_12         : out    vl_logic;
        W_53_13         : out    vl_logic;
        W_53_14         : out    vl_logic;
        W_53_15         : out    vl_logic;
        W_53_16         : out    vl_logic;
        W_53_17         : out    vl_logic;
        W_53_18         : out    vl_logic;
        W_53_19         : out    vl_logic;
        W_53_20         : out    vl_logic;
        W_53_21         : out    vl_logic;
        W_53_22         : out    vl_logic;
        W_53_23         : out    vl_logic;
        W_53_24         : out    vl_logic;
        W_53_25         : out    vl_logic;
        W_53_26         : out    vl_logic;
        W_53_27         : out    vl_logic;
        W_53_28         : out    vl_logic;
        W_53_29         : out    vl_logic;
        W_53_30         : out    vl_logic;
        W_53_31         : out    vl_logic;
        W_52_0          : out    vl_logic;
        W_52_1          : out    vl_logic;
        W_52_2          : out    vl_logic;
        W_52_3          : out    vl_logic;
        W_52_4          : out    vl_logic;
        W_52_5          : out    vl_logic;
        W_52_6          : out    vl_logic;
        W_52_7          : out    vl_logic;
        W_52_8          : out    vl_logic;
        W_52_9          : out    vl_logic;
        W_52_10         : out    vl_logic;
        W_52_11         : out    vl_logic;
        W_52_12         : out    vl_logic;
        W_52_13         : out    vl_logic;
        W_52_14         : out    vl_logic;
        W_52_15         : out    vl_logic;
        W_52_16         : out    vl_logic;
        W_52_17         : out    vl_logic;
        W_52_18         : out    vl_logic;
        W_52_19         : out    vl_logic;
        W_52_20         : out    vl_logic;
        W_52_21         : out    vl_logic;
        W_52_22         : out    vl_logic;
        W_52_23         : out    vl_logic;
        W_52_24         : out    vl_logic;
        W_52_25         : out    vl_logic;
        W_52_26         : out    vl_logic;
        W_52_27         : out    vl_logic;
        W_52_28         : out    vl_logic;
        W_52_29         : out    vl_logic;
        W_52_30         : out    vl_logic;
        W_52_31         : out    vl_logic;
        W_51_0          : out    vl_logic;
        W_51_1          : out    vl_logic;
        W_51_2          : out    vl_logic;
        W_51_3          : out    vl_logic;
        W_51_4          : out    vl_logic;
        W_51_5          : out    vl_logic;
        W_51_6          : out    vl_logic;
        W_51_7          : out    vl_logic;
        W_51_8          : out    vl_logic;
        W_51_9          : out    vl_logic;
        W_51_10         : out    vl_logic;
        W_51_11         : out    vl_logic;
        W_51_12         : out    vl_logic;
        W_51_13         : out    vl_logic;
        W_51_14         : out    vl_logic;
        W_51_15         : out    vl_logic;
        W_51_16         : out    vl_logic;
        W_51_17         : out    vl_logic;
        W_51_18         : out    vl_logic;
        W_51_19         : out    vl_logic;
        W_51_20         : out    vl_logic;
        W_51_21         : out    vl_logic;
        W_51_22         : out    vl_logic;
        W_51_23         : out    vl_logic;
        W_51_24         : out    vl_logic;
        W_51_25         : out    vl_logic;
        W_51_26         : out    vl_logic;
        W_51_27         : out    vl_logic;
        W_51_28         : out    vl_logic;
        W_51_29         : out    vl_logic;
        W_51_30         : out    vl_logic;
        W_51_31         : out    vl_logic;
        W_50_0          : out    vl_logic;
        W_50_1          : out    vl_logic;
        W_50_2          : out    vl_logic;
        W_50_3          : out    vl_logic;
        W_50_4          : out    vl_logic;
        W_50_5          : out    vl_logic;
        W_50_6          : out    vl_logic;
        W_50_7          : out    vl_logic;
        W_50_8          : out    vl_logic;
        W_50_9          : out    vl_logic;
        W_50_10         : out    vl_logic;
        W_50_11         : out    vl_logic;
        W_50_12         : out    vl_logic;
        W_50_13         : out    vl_logic;
        W_50_14         : out    vl_logic;
        W_50_15         : out    vl_logic;
        W_50_16         : out    vl_logic;
        W_50_17         : out    vl_logic;
        W_50_18         : out    vl_logic;
        W_50_19         : out    vl_logic;
        W_50_20         : out    vl_logic;
        W_50_21         : out    vl_logic;
        W_50_22         : out    vl_logic;
        W_50_23         : out    vl_logic;
        W_50_24         : out    vl_logic;
        W_50_25         : out    vl_logic;
        W_50_26         : out    vl_logic;
        W_50_27         : out    vl_logic;
        W_50_28         : out    vl_logic;
        W_50_29         : out    vl_logic;
        W_50_30         : out    vl_logic;
        W_50_31         : out    vl_logic;
        W_49_0          : out    vl_logic;
        W_49_1          : out    vl_logic;
        W_49_2          : out    vl_logic;
        W_49_3          : out    vl_logic;
        W_49_4          : out    vl_logic;
        W_49_5          : out    vl_logic;
        W_49_6          : out    vl_logic;
        W_49_7          : out    vl_logic;
        W_49_8          : out    vl_logic;
        W_49_9          : out    vl_logic;
        W_49_10         : out    vl_logic;
        W_49_11         : out    vl_logic;
        W_49_12         : out    vl_logic;
        W_49_13         : out    vl_logic;
        W_49_14         : out    vl_logic;
        W_49_15         : out    vl_logic;
        W_49_16         : out    vl_logic;
        W_49_17         : out    vl_logic;
        W_49_18         : out    vl_logic;
        W_49_19         : out    vl_logic;
        W_49_20         : out    vl_logic;
        W_49_21         : out    vl_logic;
        W_49_22         : out    vl_logic;
        W_49_23         : out    vl_logic;
        W_49_24         : out    vl_logic;
        W_49_25         : out    vl_logic;
        W_49_26         : out    vl_logic;
        W_49_27         : out    vl_logic;
        W_49_28         : out    vl_logic;
        W_49_29         : out    vl_logic;
        W_49_30         : out    vl_logic;
        W_49_31         : out    vl_logic;
        W_48_0          : out    vl_logic;
        W_48_1          : out    vl_logic;
        W_48_2          : out    vl_logic;
        W_48_3          : out    vl_logic;
        W_48_4          : out    vl_logic;
        W_48_5          : out    vl_logic;
        W_48_6          : out    vl_logic;
        W_48_7          : out    vl_logic;
        W_48_8          : out    vl_logic;
        W_48_9          : out    vl_logic;
        W_48_10         : out    vl_logic;
        W_48_11         : out    vl_logic;
        W_48_12         : out    vl_logic;
        W_48_13         : out    vl_logic;
        W_48_14         : out    vl_logic;
        W_48_15         : out    vl_logic;
        W_48_16         : out    vl_logic;
        W_48_17         : out    vl_logic;
        W_48_18         : out    vl_logic;
        W_48_19         : out    vl_logic;
        W_48_20         : out    vl_logic;
        W_48_21         : out    vl_logic;
        W_48_22         : out    vl_logic;
        W_48_23         : out    vl_logic;
        W_48_24         : out    vl_logic;
        W_48_25         : out    vl_logic;
        W_48_26         : out    vl_logic;
        W_48_27         : out    vl_logic;
        W_48_28         : out    vl_logic;
        W_48_29         : out    vl_logic;
        W_48_30         : out    vl_logic;
        W_48_31         : out    vl_logic;
        W_47_0          : out    vl_logic;
        W_47_1          : out    vl_logic;
        W_47_2          : out    vl_logic;
        W_47_3          : out    vl_logic;
        W_47_4          : out    vl_logic;
        W_47_5          : out    vl_logic;
        W_47_6          : out    vl_logic;
        W_47_7          : out    vl_logic;
        W_47_8          : out    vl_logic;
        W_47_9          : out    vl_logic;
        W_47_10         : out    vl_logic;
        W_47_11         : out    vl_logic;
        W_47_12         : out    vl_logic;
        W_47_13         : out    vl_logic;
        W_47_14         : out    vl_logic;
        W_47_15         : out    vl_logic;
        W_47_16         : out    vl_logic;
        W_47_17         : out    vl_logic;
        W_47_18         : out    vl_logic;
        W_47_19         : out    vl_logic;
        W_47_20         : out    vl_logic;
        W_47_21         : out    vl_logic;
        W_47_22         : out    vl_logic;
        W_47_23         : out    vl_logic;
        W_47_24         : out    vl_logic;
        W_47_25         : out    vl_logic;
        W_47_26         : out    vl_logic;
        W_47_27         : out    vl_logic;
        W_47_28         : out    vl_logic;
        W_47_29         : out    vl_logic;
        W_47_30         : out    vl_logic;
        W_47_31         : out    vl_logic;
        W_46_0          : out    vl_logic;
        W_46_1          : out    vl_logic;
        W_46_2          : out    vl_logic;
        W_46_3          : out    vl_logic;
        W_46_4          : out    vl_logic;
        W_46_5          : out    vl_logic;
        W_46_6          : out    vl_logic;
        W_46_7          : out    vl_logic;
        W_46_8          : out    vl_logic;
        W_46_9          : out    vl_logic;
        W_46_10         : out    vl_logic;
        W_46_11         : out    vl_logic;
        W_46_12         : out    vl_logic;
        W_46_13         : out    vl_logic;
        W_46_14         : out    vl_logic;
        W_46_15         : out    vl_logic;
        W_46_16         : out    vl_logic;
        W_46_17         : out    vl_logic;
        W_46_18         : out    vl_logic;
        W_46_19         : out    vl_logic;
        W_46_20         : out    vl_logic;
        W_46_21         : out    vl_logic;
        W_46_22         : out    vl_logic;
        W_46_23         : out    vl_logic;
        W_46_24         : out    vl_logic;
        W_46_25         : out    vl_logic;
        W_46_26         : out    vl_logic;
        W_46_27         : out    vl_logic;
        W_46_28         : out    vl_logic;
        W_46_29         : out    vl_logic;
        W_46_30         : out    vl_logic;
        W_46_31         : out    vl_logic;
        W_45_0          : out    vl_logic;
        W_45_1          : out    vl_logic;
        W_45_2          : out    vl_logic;
        W_45_3          : out    vl_logic;
        W_45_4          : out    vl_logic;
        W_45_5          : out    vl_logic;
        W_45_6          : out    vl_logic;
        W_45_7          : out    vl_logic;
        W_45_8          : out    vl_logic;
        W_45_9          : out    vl_logic;
        W_45_10         : out    vl_logic;
        W_45_11         : out    vl_logic;
        W_45_12         : out    vl_logic;
        W_45_13         : out    vl_logic;
        W_45_14         : out    vl_logic;
        W_45_15         : out    vl_logic;
        W_45_16         : out    vl_logic;
        W_45_17         : out    vl_logic;
        W_45_18         : out    vl_logic;
        W_45_19         : out    vl_logic;
        W_45_20         : out    vl_logic;
        W_45_21         : out    vl_logic;
        W_45_22         : out    vl_logic;
        W_45_23         : out    vl_logic;
        W_45_24         : out    vl_logic;
        W_45_25         : out    vl_logic;
        W_45_26         : out    vl_logic;
        W_45_27         : out    vl_logic;
        W_45_28         : out    vl_logic;
        W_45_29         : out    vl_logic;
        W_45_30         : out    vl_logic;
        W_45_31         : out    vl_logic;
        W_44_0          : out    vl_logic;
        W_44_1          : out    vl_logic;
        W_44_2          : out    vl_logic;
        W_44_3          : out    vl_logic;
        W_44_4          : out    vl_logic;
        W_44_5          : out    vl_logic;
        W_44_6          : out    vl_logic;
        W_44_7          : out    vl_logic;
        W_44_8          : out    vl_logic;
        W_44_9          : out    vl_logic;
        W_44_10         : out    vl_logic;
        W_44_11         : out    vl_logic;
        W_44_12         : out    vl_logic;
        W_44_13         : out    vl_logic;
        W_44_14         : out    vl_logic;
        W_44_15         : out    vl_logic;
        W_44_16         : out    vl_logic;
        W_44_17         : out    vl_logic;
        W_44_18         : out    vl_logic;
        W_44_19         : out    vl_logic;
        W_44_20         : out    vl_logic;
        W_44_21         : out    vl_logic;
        W_44_22         : out    vl_logic;
        W_44_23         : out    vl_logic;
        W_44_24         : out    vl_logic;
        W_44_25         : out    vl_logic;
        W_44_26         : out    vl_logic;
        W_44_27         : out    vl_logic;
        W_44_28         : out    vl_logic;
        W_44_29         : out    vl_logic;
        W_44_30         : out    vl_logic;
        W_44_31         : out    vl_logic;
        W_43_0          : out    vl_logic;
        W_43_1          : out    vl_logic;
        W_43_2          : out    vl_logic;
        W_43_3          : out    vl_logic;
        W_43_4          : out    vl_logic;
        W_43_5          : out    vl_logic;
        W_43_6          : out    vl_logic;
        W_43_7          : out    vl_logic;
        W_43_8          : out    vl_logic;
        W_43_9          : out    vl_logic;
        W_43_10         : out    vl_logic;
        W_43_11         : out    vl_logic;
        W_43_12         : out    vl_logic;
        W_43_13         : out    vl_logic;
        W_43_14         : out    vl_logic;
        W_43_15         : out    vl_logic;
        W_43_16         : out    vl_logic;
        W_43_17         : out    vl_logic;
        W_43_18         : out    vl_logic;
        W_43_19         : out    vl_logic;
        W_43_20         : out    vl_logic;
        W_43_21         : out    vl_logic;
        W_43_22         : out    vl_logic;
        W_43_23         : out    vl_logic;
        W_43_24         : out    vl_logic;
        W_43_25         : out    vl_logic;
        W_43_26         : out    vl_logic;
        W_43_27         : out    vl_logic;
        W_43_28         : out    vl_logic;
        W_43_29         : out    vl_logic;
        W_43_30         : out    vl_logic;
        W_43_31         : out    vl_logic;
        W_42_0          : out    vl_logic;
        W_42_1          : out    vl_logic;
        W_42_2          : out    vl_logic;
        W_42_3          : out    vl_logic;
        W_42_4          : out    vl_logic;
        W_42_5          : out    vl_logic;
        W_42_6          : out    vl_logic;
        W_42_7          : out    vl_logic;
        W_42_8          : out    vl_logic;
        W_42_9          : out    vl_logic;
        W_42_10         : out    vl_logic;
        W_42_11         : out    vl_logic;
        W_42_12         : out    vl_logic;
        W_42_13         : out    vl_logic;
        W_42_14         : out    vl_logic;
        W_42_15         : out    vl_logic;
        W_42_16         : out    vl_logic;
        W_42_17         : out    vl_logic;
        W_42_18         : out    vl_logic;
        W_42_19         : out    vl_logic;
        W_42_20         : out    vl_logic;
        W_42_21         : out    vl_logic;
        W_42_22         : out    vl_logic;
        W_42_23         : out    vl_logic;
        W_42_24         : out    vl_logic;
        W_42_25         : out    vl_logic;
        W_42_26         : out    vl_logic;
        W_42_27         : out    vl_logic;
        W_42_28         : out    vl_logic;
        W_42_29         : out    vl_logic;
        W_42_30         : out    vl_logic;
        W_42_31         : out    vl_logic;
        W_41_0          : out    vl_logic;
        W_41_1          : out    vl_logic;
        W_41_2          : out    vl_logic;
        W_41_3          : out    vl_logic;
        W_41_4          : out    vl_logic;
        W_41_5          : out    vl_logic;
        W_41_6          : out    vl_logic;
        W_41_7          : out    vl_logic;
        W_41_8          : out    vl_logic;
        W_41_9          : out    vl_logic;
        W_41_10         : out    vl_logic;
        W_41_11         : out    vl_logic;
        W_41_12         : out    vl_logic;
        W_41_13         : out    vl_logic;
        W_41_14         : out    vl_logic;
        W_41_15         : out    vl_logic;
        W_41_16         : out    vl_logic;
        W_41_17         : out    vl_logic;
        W_41_18         : out    vl_logic;
        W_41_19         : out    vl_logic;
        W_41_20         : out    vl_logic;
        W_41_21         : out    vl_logic;
        W_41_22         : out    vl_logic;
        W_41_23         : out    vl_logic;
        W_41_24         : out    vl_logic;
        W_41_25         : out    vl_logic;
        W_41_26         : out    vl_logic;
        W_41_27         : out    vl_logic;
        W_41_28         : out    vl_logic;
        W_41_29         : out    vl_logic;
        W_41_30         : out    vl_logic;
        W_41_31         : out    vl_logic;
        W_40_0          : out    vl_logic;
        W_40_1          : out    vl_logic;
        W_40_2          : out    vl_logic;
        W_40_3          : out    vl_logic;
        W_40_4          : out    vl_logic;
        W_40_5          : out    vl_logic;
        W_40_6          : out    vl_logic;
        W_40_7          : out    vl_logic;
        W_40_8          : out    vl_logic;
        W_40_9          : out    vl_logic;
        W_40_10         : out    vl_logic;
        W_40_11         : out    vl_logic;
        W_40_12         : out    vl_logic;
        W_40_13         : out    vl_logic;
        W_40_14         : out    vl_logic;
        W_40_15         : out    vl_logic;
        W_40_16         : out    vl_logic;
        W_40_17         : out    vl_logic;
        W_40_18         : out    vl_logic;
        W_40_19         : out    vl_logic;
        W_40_20         : out    vl_logic;
        W_40_21         : out    vl_logic;
        W_40_22         : out    vl_logic;
        W_40_23         : out    vl_logic;
        W_40_24         : out    vl_logic;
        W_40_25         : out    vl_logic;
        W_40_26         : out    vl_logic;
        W_40_27         : out    vl_logic;
        W_40_28         : out    vl_logic;
        W_40_29         : out    vl_logic;
        W_40_30         : out    vl_logic;
        W_40_31         : out    vl_logic;
        W_39_0          : out    vl_logic;
        W_39_1          : out    vl_logic;
        W_39_2          : out    vl_logic;
        W_39_3          : out    vl_logic;
        W_39_4          : out    vl_logic;
        W_39_5          : out    vl_logic;
        W_39_6          : out    vl_logic;
        W_39_7          : out    vl_logic;
        W_39_8          : out    vl_logic;
        W_39_9          : out    vl_logic;
        W_39_10         : out    vl_logic;
        W_39_11         : out    vl_logic;
        W_39_12         : out    vl_logic;
        W_39_13         : out    vl_logic;
        W_39_14         : out    vl_logic;
        W_39_15         : out    vl_logic;
        W_39_16         : out    vl_logic;
        W_39_17         : out    vl_logic;
        W_39_18         : out    vl_logic;
        W_39_19         : out    vl_logic;
        W_39_20         : out    vl_logic;
        W_39_21         : out    vl_logic;
        W_39_22         : out    vl_logic;
        W_39_23         : out    vl_logic;
        W_39_24         : out    vl_logic;
        W_39_25         : out    vl_logic;
        W_39_26         : out    vl_logic;
        W_39_27         : out    vl_logic;
        W_39_28         : out    vl_logic;
        W_39_29         : out    vl_logic;
        W_39_30         : out    vl_logic;
        W_39_31         : out    vl_logic;
        W_38_0          : out    vl_logic;
        W_38_1          : out    vl_logic;
        W_38_2          : out    vl_logic;
        W_38_3          : out    vl_logic;
        W_38_4          : out    vl_logic;
        W_38_5          : out    vl_logic;
        W_38_6          : out    vl_logic;
        W_38_7          : out    vl_logic;
        W_38_8          : out    vl_logic;
        W_38_9          : out    vl_logic;
        W_38_10         : out    vl_logic;
        W_38_11         : out    vl_logic;
        W_38_12         : out    vl_logic;
        W_38_13         : out    vl_logic;
        W_38_14         : out    vl_logic;
        W_38_15         : out    vl_logic;
        W_38_16         : out    vl_logic;
        W_38_17         : out    vl_logic;
        W_38_18         : out    vl_logic;
        W_38_19         : out    vl_logic;
        W_38_20         : out    vl_logic;
        W_38_21         : out    vl_logic;
        W_38_22         : out    vl_logic;
        W_38_23         : out    vl_logic;
        W_38_24         : out    vl_logic;
        W_38_25         : out    vl_logic;
        W_38_26         : out    vl_logic;
        W_38_27         : out    vl_logic;
        W_38_28         : out    vl_logic;
        W_38_29         : out    vl_logic;
        W_38_30         : out    vl_logic;
        W_38_31         : out    vl_logic;
        W_37_0          : out    vl_logic;
        W_37_1          : out    vl_logic;
        W_37_2          : out    vl_logic;
        W_37_3          : out    vl_logic;
        W_37_4          : out    vl_logic;
        W_37_5          : out    vl_logic;
        W_37_6          : out    vl_logic;
        W_37_7          : out    vl_logic;
        W_37_8          : out    vl_logic;
        W_37_9          : out    vl_logic;
        W_37_10         : out    vl_logic;
        W_37_11         : out    vl_logic;
        W_37_12         : out    vl_logic;
        W_37_13         : out    vl_logic;
        W_37_14         : out    vl_logic;
        W_37_15         : out    vl_logic;
        W_37_16         : out    vl_logic;
        W_37_17         : out    vl_logic;
        W_37_18         : out    vl_logic;
        W_37_19         : out    vl_logic;
        W_37_20         : out    vl_logic;
        W_37_21         : out    vl_logic;
        W_37_22         : out    vl_logic;
        W_37_23         : out    vl_logic;
        W_37_24         : out    vl_logic;
        W_37_25         : out    vl_logic;
        W_37_26         : out    vl_logic;
        W_37_27         : out    vl_logic;
        W_37_28         : out    vl_logic;
        W_37_29         : out    vl_logic;
        W_37_30         : out    vl_logic;
        W_37_31         : out    vl_logic;
        W_36_0          : out    vl_logic;
        W_36_1          : out    vl_logic;
        W_36_2          : out    vl_logic;
        W_36_3          : out    vl_logic;
        W_36_4          : out    vl_logic;
        W_36_5          : out    vl_logic;
        W_36_6          : out    vl_logic;
        W_36_7          : out    vl_logic;
        W_36_8          : out    vl_logic;
        W_36_9          : out    vl_logic;
        W_36_10         : out    vl_logic;
        W_36_11         : out    vl_logic;
        W_36_12         : out    vl_logic;
        W_36_13         : out    vl_logic;
        W_36_14         : out    vl_logic;
        W_36_15         : out    vl_logic;
        W_36_16         : out    vl_logic;
        W_36_17         : out    vl_logic;
        W_36_18         : out    vl_logic;
        W_36_19         : out    vl_logic;
        W_36_20         : out    vl_logic;
        W_36_21         : out    vl_logic;
        W_36_22         : out    vl_logic;
        W_36_23         : out    vl_logic;
        W_36_24         : out    vl_logic;
        W_36_25         : out    vl_logic;
        W_36_26         : out    vl_logic;
        W_36_27         : out    vl_logic;
        W_36_28         : out    vl_logic;
        W_36_29         : out    vl_logic;
        W_36_30         : out    vl_logic;
        W_36_31         : out    vl_logic;
        W_35_0          : out    vl_logic;
        W_35_1          : out    vl_logic;
        W_35_2          : out    vl_logic;
        W_35_3          : out    vl_logic;
        W_35_4          : out    vl_logic;
        W_35_5          : out    vl_logic;
        W_35_6          : out    vl_logic;
        W_35_7          : out    vl_logic;
        W_35_8          : out    vl_logic;
        W_35_9          : out    vl_logic;
        W_35_10         : out    vl_logic;
        W_35_11         : out    vl_logic;
        W_35_12         : out    vl_logic;
        W_35_13         : out    vl_logic;
        W_35_14         : out    vl_logic;
        W_35_15         : out    vl_logic;
        W_35_16         : out    vl_logic;
        W_35_17         : out    vl_logic;
        W_35_18         : out    vl_logic;
        W_35_19         : out    vl_logic;
        W_35_20         : out    vl_logic;
        W_35_21         : out    vl_logic;
        W_35_22         : out    vl_logic;
        W_35_23         : out    vl_logic;
        W_35_24         : out    vl_logic;
        W_35_25         : out    vl_logic;
        W_35_26         : out    vl_logic;
        W_35_27         : out    vl_logic;
        W_35_28         : out    vl_logic;
        W_35_29         : out    vl_logic;
        W_35_30         : out    vl_logic;
        W_35_31         : out    vl_logic;
        W_34_0          : out    vl_logic;
        W_34_1          : out    vl_logic;
        W_34_2          : out    vl_logic;
        W_34_3          : out    vl_logic;
        W_34_4          : out    vl_logic;
        W_34_5          : out    vl_logic;
        W_34_6          : out    vl_logic;
        W_34_7          : out    vl_logic;
        W_34_8          : out    vl_logic;
        W_34_9          : out    vl_logic;
        W_34_10         : out    vl_logic;
        W_34_11         : out    vl_logic;
        W_34_12         : out    vl_logic;
        W_34_13         : out    vl_logic;
        W_34_14         : out    vl_logic;
        W_34_15         : out    vl_logic;
        W_34_16         : out    vl_logic;
        W_34_17         : out    vl_logic;
        W_34_18         : out    vl_logic;
        W_34_19         : out    vl_logic;
        W_34_20         : out    vl_logic;
        W_34_21         : out    vl_logic;
        W_34_22         : out    vl_logic;
        W_34_23         : out    vl_logic;
        W_34_24         : out    vl_logic;
        W_34_25         : out    vl_logic;
        W_34_26         : out    vl_logic;
        W_34_27         : out    vl_logic;
        W_34_28         : out    vl_logic;
        W_34_29         : out    vl_logic;
        W_34_30         : out    vl_logic;
        W_34_31         : out    vl_logic;
        W_33_0          : out    vl_logic;
        W_33_1          : out    vl_logic;
        W_33_2          : out    vl_logic;
        W_33_3          : out    vl_logic;
        W_33_4          : out    vl_logic;
        W_33_5          : out    vl_logic;
        W_33_6          : out    vl_logic;
        W_33_7          : out    vl_logic;
        W_33_8          : out    vl_logic;
        W_33_9          : out    vl_logic;
        W_33_10         : out    vl_logic;
        W_33_11         : out    vl_logic;
        W_33_12         : out    vl_logic;
        W_33_13         : out    vl_logic;
        W_33_14         : out    vl_logic;
        W_33_15         : out    vl_logic;
        W_33_16         : out    vl_logic;
        W_33_17         : out    vl_logic;
        W_33_18         : out    vl_logic;
        W_33_19         : out    vl_logic;
        W_33_20         : out    vl_logic;
        W_33_21         : out    vl_logic;
        W_33_22         : out    vl_logic;
        W_33_23         : out    vl_logic;
        W_33_24         : out    vl_logic;
        W_33_25         : out    vl_logic;
        W_33_26         : out    vl_logic;
        W_33_27         : out    vl_logic;
        W_33_28         : out    vl_logic;
        W_33_29         : out    vl_logic;
        W_33_30         : out    vl_logic;
        W_33_31         : out    vl_logic;
        W_32_0          : out    vl_logic;
        W_32_1          : out    vl_logic;
        W_32_2          : out    vl_logic;
        W_32_3          : out    vl_logic;
        W_32_4          : out    vl_logic;
        W_32_5          : out    vl_logic;
        W_32_6          : out    vl_logic;
        W_32_7          : out    vl_logic;
        W_32_8          : out    vl_logic;
        W_32_9          : out    vl_logic;
        W_32_10         : out    vl_logic;
        W_32_11         : out    vl_logic;
        W_32_12         : out    vl_logic;
        W_32_13         : out    vl_logic;
        W_32_14         : out    vl_logic;
        W_32_15         : out    vl_logic;
        W_32_16         : out    vl_logic;
        W_32_17         : out    vl_logic;
        W_32_18         : out    vl_logic;
        W_32_19         : out    vl_logic;
        W_32_20         : out    vl_logic;
        W_32_21         : out    vl_logic;
        W_32_22         : out    vl_logic;
        W_32_23         : out    vl_logic;
        W_32_24         : out    vl_logic;
        W_32_25         : out    vl_logic;
        W_32_26         : out    vl_logic;
        W_32_27         : out    vl_logic;
        W_32_28         : out    vl_logic;
        W_32_29         : out    vl_logic;
        W_32_30         : out    vl_logic;
        W_32_31         : out    vl_logic;
        W_31_0          : out    vl_logic;
        W_31_1          : out    vl_logic;
        W_31_2          : out    vl_logic;
        W_31_3          : out    vl_logic;
        W_31_4          : out    vl_logic;
        W_31_5          : out    vl_logic;
        W_31_6          : out    vl_logic;
        W_31_7          : out    vl_logic;
        W_31_8          : out    vl_logic;
        W_31_9          : out    vl_logic;
        W_31_10         : out    vl_logic;
        W_31_11         : out    vl_logic;
        W_31_12         : out    vl_logic;
        W_31_13         : out    vl_logic;
        W_31_14         : out    vl_logic;
        W_31_15         : out    vl_logic;
        W_31_16         : out    vl_logic;
        W_31_17         : out    vl_logic;
        W_31_18         : out    vl_logic;
        W_31_19         : out    vl_logic;
        W_31_20         : out    vl_logic;
        W_31_21         : out    vl_logic;
        W_31_22         : out    vl_logic;
        W_31_23         : out    vl_logic;
        W_31_24         : out    vl_logic;
        W_31_25         : out    vl_logic;
        W_31_26         : out    vl_logic;
        W_31_27         : out    vl_logic;
        W_31_28         : out    vl_logic;
        W_31_29         : out    vl_logic;
        W_31_30         : out    vl_logic;
        W_31_31         : out    vl_logic;
        W_30_0          : out    vl_logic;
        W_30_1          : out    vl_logic;
        W_30_2          : out    vl_logic;
        W_30_3          : out    vl_logic;
        W_30_4          : out    vl_logic;
        W_30_5          : out    vl_logic;
        W_30_6          : out    vl_logic;
        W_30_7          : out    vl_logic;
        W_30_8          : out    vl_logic;
        W_30_9          : out    vl_logic;
        W_30_10         : out    vl_logic;
        W_30_11         : out    vl_logic;
        W_30_12         : out    vl_logic;
        W_30_13         : out    vl_logic;
        W_30_14         : out    vl_logic;
        W_30_15         : out    vl_logic;
        W_30_16         : out    vl_logic;
        W_30_17         : out    vl_logic;
        W_30_18         : out    vl_logic;
        W_30_19         : out    vl_logic;
        W_30_20         : out    vl_logic;
        W_30_21         : out    vl_logic;
        W_30_22         : out    vl_logic;
        W_30_23         : out    vl_logic;
        W_30_24         : out    vl_logic;
        W_30_25         : out    vl_logic;
        W_30_26         : out    vl_logic;
        W_30_27         : out    vl_logic;
        W_30_28         : out    vl_logic;
        W_30_29         : out    vl_logic;
        W_30_30         : out    vl_logic;
        W_30_31         : out    vl_logic;
        W_29_0          : out    vl_logic;
        W_29_1          : out    vl_logic;
        W_29_2          : out    vl_logic;
        W_29_3          : out    vl_logic;
        W_29_4          : out    vl_logic;
        W_29_5          : out    vl_logic;
        W_29_6          : out    vl_logic;
        W_29_7          : out    vl_logic;
        W_29_8          : out    vl_logic;
        W_29_9          : out    vl_logic;
        W_29_10         : out    vl_logic;
        W_29_11         : out    vl_logic;
        W_29_12         : out    vl_logic;
        W_29_13         : out    vl_logic;
        W_29_14         : out    vl_logic;
        W_29_15         : out    vl_logic;
        W_29_16         : out    vl_logic;
        W_29_17         : out    vl_logic;
        W_29_18         : out    vl_logic;
        W_29_19         : out    vl_logic;
        W_29_20         : out    vl_logic;
        W_29_21         : out    vl_logic;
        W_29_22         : out    vl_logic;
        W_29_23         : out    vl_logic;
        W_29_24         : out    vl_logic;
        W_29_25         : out    vl_logic;
        W_29_26         : out    vl_logic;
        W_29_27         : out    vl_logic;
        W_29_28         : out    vl_logic;
        W_29_29         : out    vl_logic;
        W_29_30         : out    vl_logic;
        W_29_31         : out    vl_logic;
        W_28_0          : out    vl_logic;
        W_28_1          : out    vl_logic;
        W_28_2          : out    vl_logic;
        W_28_3          : out    vl_logic;
        W_28_4          : out    vl_logic;
        W_28_5          : out    vl_logic;
        W_28_6          : out    vl_logic;
        W_28_7          : out    vl_logic;
        W_28_8          : out    vl_logic;
        W_28_9          : out    vl_logic;
        W_28_10         : out    vl_logic;
        W_28_11         : out    vl_logic;
        W_28_12         : out    vl_logic;
        W_28_13         : out    vl_logic;
        W_28_14         : out    vl_logic;
        W_28_15         : out    vl_logic;
        W_28_16         : out    vl_logic;
        W_28_17         : out    vl_logic;
        W_28_18         : out    vl_logic;
        W_28_19         : out    vl_logic;
        W_28_20         : out    vl_logic;
        W_28_21         : out    vl_logic;
        W_28_22         : out    vl_logic;
        W_28_23         : out    vl_logic;
        W_28_24         : out    vl_logic;
        W_28_25         : out    vl_logic;
        W_28_26         : out    vl_logic;
        W_28_27         : out    vl_logic;
        W_28_28         : out    vl_logic;
        W_28_29         : out    vl_logic;
        W_28_30         : out    vl_logic;
        W_28_31         : out    vl_logic;
        W_27_0          : out    vl_logic;
        W_27_1          : out    vl_logic;
        W_27_2          : out    vl_logic;
        W_27_3          : out    vl_logic;
        W_27_4          : out    vl_logic;
        W_27_5          : out    vl_logic;
        W_27_6          : out    vl_logic;
        W_27_7          : out    vl_logic;
        W_27_8          : out    vl_logic;
        W_27_9          : out    vl_logic;
        W_27_10         : out    vl_logic;
        W_27_11         : out    vl_logic;
        W_27_12         : out    vl_logic;
        W_27_13         : out    vl_logic;
        W_27_14         : out    vl_logic;
        W_27_15         : out    vl_logic;
        W_27_16         : out    vl_logic;
        W_27_17         : out    vl_logic;
        W_27_18         : out    vl_logic;
        W_27_19         : out    vl_logic;
        W_27_20         : out    vl_logic;
        W_27_21         : out    vl_logic;
        W_27_22         : out    vl_logic;
        W_27_23         : out    vl_logic;
        W_27_24         : out    vl_logic;
        W_27_25         : out    vl_logic;
        W_27_26         : out    vl_logic;
        W_27_27         : out    vl_logic;
        W_27_28         : out    vl_logic;
        W_27_29         : out    vl_logic;
        W_27_30         : out    vl_logic;
        W_27_31         : out    vl_logic;
        W_26_0          : out    vl_logic;
        W_26_1          : out    vl_logic;
        W_26_2          : out    vl_logic;
        W_26_3          : out    vl_logic;
        W_26_4          : out    vl_logic;
        W_26_5          : out    vl_logic;
        W_26_6          : out    vl_logic;
        W_26_7          : out    vl_logic;
        W_26_8          : out    vl_logic;
        W_26_9          : out    vl_logic;
        W_26_10         : out    vl_logic;
        W_26_11         : out    vl_logic;
        W_26_12         : out    vl_logic;
        W_26_13         : out    vl_logic;
        W_26_14         : out    vl_logic;
        W_26_15         : out    vl_logic;
        W_26_16         : out    vl_logic;
        W_26_17         : out    vl_logic;
        W_26_18         : out    vl_logic;
        W_26_19         : out    vl_logic;
        W_26_20         : out    vl_logic;
        W_26_21         : out    vl_logic;
        W_26_22         : out    vl_logic;
        W_26_23         : out    vl_logic;
        W_26_24         : out    vl_logic;
        W_26_25         : out    vl_logic;
        W_26_26         : out    vl_logic;
        W_26_27         : out    vl_logic;
        W_26_28         : out    vl_logic;
        W_26_29         : out    vl_logic;
        W_26_30         : out    vl_logic;
        W_26_31         : out    vl_logic;
        W_25_0          : out    vl_logic;
        W_25_1          : out    vl_logic;
        W_25_2          : out    vl_logic;
        W_25_3          : out    vl_logic;
        W_25_4          : out    vl_logic;
        W_25_5          : out    vl_logic;
        W_25_6          : out    vl_logic;
        W_25_7          : out    vl_logic;
        W_25_8          : out    vl_logic;
        W_25_9          : out    vl_logic;
        W_25_10         : out    vl_logic;
        W_25_11         : out    vl_logic;
        W_25_12         : out    vl_logic;
        W_25_13         : out    vl_logic;
        W_25_14         : out    vl_logic;
        W_25_15         : out    vl_logic;
        W_25_16         : out    vl_logic;
        W_25_17         : out    vl_logic;
        W_25_18         : out    vl_logic;
        W_25_19         : out    vl_logic;
        W_25_20         : out    vl_logic;
        W_25_21         : out    vl_logic;
        W_25_22         : out    vl_logic;
        W_25_23         : out    vl_logic;
        W_25_24         : out    vl_logic;
        W_25_25         : out    vl_logic;
        W_25_26         : out    vl_logic;
        W_25_27         : out    vl_logic;
        W_25_28         : out    vl_logic;
        W_25_29         : out    vl_logic;
        W_25_30         : out    vl_logic;
        W_25_31         : out    vl_logic;
        W_24_0          : out    vl_logic;
        W_24_1          : out    vl_logic;
        W_24_2          : out    vl_logic;
        W_24_3          : out    vl_logic;
        W_24_4          : out    vl_logic;
        W_24_5          : out    vl_logic;
        W_24_6          : out    vl_logic;
        W_24_7          : out    vl_logic;
        W_24_8          : out    vl_logic;
        W_24_9          : out    vl_logic;
        W_24_10         : out    vl_logic;
        W_24_11         : out    vl_logic;
        W_24_12         : out    vl_logic;
        W_24_13         : out    vl_logic;
        W_24_14         : out    vl_logic;
        W_24_15         : out    vl_logic;
        W_24_16         : out    vl_logic;
        W_24_17         : out    vl_logic;
        W_24_18         : out    vl_logic;
        W_24_19         : out    vl_logic;
        W_24_20         : out    vl_logic;
        W_24_21         : out    vl_logic;
        W_24_22         : out    vl_logic;
        W_24_23         : out    vl_logic;
        W_24_24         : out    vl_logic;
        W_24_25         : out    vl_logic;
        W_24_26         : out    vl_logic;
        W_24_27         : out    vl_logic;
        W_24_28         : out    vl_logic;
        W_24_29         : out    vl_logic;
        W_24_30         : out    vl_logic;
        W_24_31         : out    vl_logic;
        W_23_0          : out    vl_logic;
        W_23_1          : out    vl_logic;
        W_23_2          : out    vl_logic;
        W_23_3          : out    vl_logic;
        W_23_4          : out    vl_logic;
        W_23_5          : out    vl_logic;
        W_23_6          : out    vl_logic;
        W_23_7          : out    vl_logic;
        W_23_8          : out    vl_logic;
        W_23_9          : out    vl_logic;
        W_23_10         : out    vl_logic;
        W_23_11         : out    vl_logic;
        W_23_12         : out    vl_logic;
        W_23_13         : out    vl_logic;
        W_23_14         : out    vl_logic;
        W_23_15         : out    vl_logic;
        W_23_16         : out    vl_logic;
        W_23_17         : out    vl_logic;
        W_23_18         : out    vl_logic;
        W_23_19         : out    vl_logic;
        W_23_20         : out    vl_logic;
        W_23_21         : out    vl_logic;
        W_23_22         : out    vl_logic;
        W_23_23         : out    vl_logic;
        W_23_24         : out    vl_logic;
        W_23_25         : out    vl_logic;
        W_23_26         : out    vl_logic;
        W_23_27         : out    vl_logic;
        W_23_28         : out    vl_logic;
        W_23_29         : out    vl_logic;
        W_23_30         : out    vl_logic;
        W_23_31         : out    vl_logic;
        W_22_0          : out    vl_logic;
        W_22_1          : out    vl_logic;
        W_22_2          : out    vl_logic;
        W_22_3          : out    vl_logic;
        W_22_4          : out    vl_logic;
        W_22_5          : out    vl_logic;
        W_22_6          : out    vl_logic;
        W_22_7          : out    vl_logic;
        W_22_8          : out    vl_logic;
        W_22_9          : out    vl_logic;
        W_22_10         : out    vl_logic;
        W_22_11         : out    vl_logic;
        W_22_12         : out    vl_logic;
        W_22_13         : out    vl_logic;
        W_22_14         : out    vl_logic;
        W_22_15         : out    vl_logic;
        W_22_16         : out    vl_logic;
        W_22_17         : out    vl_logic;
        W_22_18         : out    vl_logic;
        W_22_19         : out    vl_logic;
        W_22_20         : out    vl_logic;
        W_22_21         : out    vl_logic;
        W_22_22         : out    vl_logic;
        W_22_23         : out    vl_logic;
        W_22_24         : out    vl_logic;
        W_22_25         : out    vl_logic;
        W_22_26         : out    vl_logic;
        W_22_27         : out    vl_logic;
        W_22_28         : out    vl_logic;
        W_22_29         : out    vl_logic;
        W_22_30         : out    vl_logic;
        W_22_31         : out    vl_logic;
        W_21_0          : out    vl_logic;
        W_21_1          : out    vl_logic;
        W_21_2          : out    vl_logic;
        W_21_3          : out    vl_logic;
        W_21_4          : out    vl_logic;
        W_21_5          : out    vl_logic;
        W_21_6          : out    vl_logic;
        W_21_7          : out    vl_logic;
        W_21_8          : out    vl_logic;
        W_21_9          : out    vl_logic;
        W_21_10         : out    vl_logic;
        W_21_11         : out    vl_logic;
        W_21_12         : out    vl_logic;
        W_21_13         : out    vl_logic;
        W_21_14         : out    vl_logic;
        W_21_15         : out    vl_logic;
        W_21_16         : out    vl_logic;
        W_21_17         : out    vl_logic;
        W_21_18         : out    vl_logic;
        W_21_19         : out    vl_logic;
        W_21_20         : out    vl_logic;
        W_21_21         : out    vl_logic;
        W_21_22         : out    vl_logic;
        W_21_23         : out    vl_logic;
        W_21_24         : out    vl_logic;
        W_21_25         : out    vl_logic;
        W_21_26         : out    vl_logic;
        W_21_27         : out    vl_logic;
        W_21_28         : out    vl_logic;
        W_21_29         : out    vl_logic;
        W_21_30         : out    vl_logic;
        W_21_31         : out    vl_logic;
        W_20_0          : out    vl_logic;
        W_20_1          : out    vl_logic;
        W_20_2          : out    vl_logic;
        W_20_3          : out    vl_logic;
        W_20_4          : out    vl_logic;
        W_20_5          : out    vl_logic;
        W_20_6          : out    vl_logic;
        W_20_7          : out    vl_logic;
        W_20_8          : out    vl_logic;
        W_20_9          : out    vl_logic;
        W_20_10         : out    vl_logic;
        W_20_11         : out    vl_logic;
        W_20_12         : out    vl_logic;
        W_20_13         : out    vl_logic;
        W_20_14         : out    vl_logic;
        W_20_15         : out    vl_logic;
        W_20_16         : out    vl_logic;
        W_20_17         : out    vl_logic;
        W_20_18         : out    vl_logic;
        W_20_19         : out    vl_logic;
        W_20_20         : out    vl_logic;
        W_20_21         : out    vl_logic;
        W_20_22         : out    vl_logic;
        W_20_23         : out    vl_logic;
        W_20_24         : out    vl_logic;
        W_20_25         : out    vl_logic;
        W_20_26         : out    vl_logic;
        W_20_27         : out    vl_logic;
        W_20_28         : out    vl_logic;
        W_20_29         : out    vl_logic;
        W_20_30         : out    vl_logic;
        W_20_31         : out    vl_logic;
        W_19_0          : out    vl_logic;
        W_19_1          : out    vl_logic;
        W_19_2          : out    vl_logic;
        W_19_3          : out    vl_logic;
        W_19_4          : out    vl_logic;
        W_19_5          : out    vl_logic;
        W_19_6          : out    vl_logic;
        W_19_7          : out    vl_logic;
        W_19_8          : out    vl_logic;
        W_19_9          : out    vl_logic;
        W_19_10         : out    vl_logic;
        W_19_11         : out    vl_logic;
        W_19_12         : out    vl_logic;
        W_19_13         : out    vl_logic;
        W_19_14         : out    vl_logic;
        W_19_15         : out    vl_logic;
        W_19_16         : out    vl_logic;
        W_19_17         : out    vl_logic;
        W_19_18         : out    vl_logic;
        W_19_19         : out    vl_logic;
        W_19_20         : out    vl_logic;
        W_19_21         : out    vl_logic;
        W_19_22         : out    vl_logic;
        W_19_23         : out    vl_logic;
        W_19_24         : out    vl_logic;
        W_19_25         : out    vl_logic;
        W_19_26         : out    vl_logic;
        W_19_27         : out    vl_logic;
        W_19_28         : out    vl_logic;
        W_19_29         : out    vl_logic;
        W_19_30         : out    vl_logic;
        W_19_31         : out    vl_logic;
        W_18_0          : out    vl_logic;
        W_18_1          : out    vl_logic;
        W_18_2          : out    vl_logic;
        W_18_3          : out    vl_logic;
        W_18_4          : out    vl_logic;
        W_18_5          : out    vl_logic;
        W_18_6          : out    vl_logic;
        W_18_7          : out    vl_logic;
        W_18_8          : out    vl_logic;
        W_18_9          : out    vl_logic;
        W_18_10         : out    vl_logic;
        W_18_11         : out    vl_logic;
        W_18_12         : out    vl_logic;
        W_18_13         : out    vl_logic;
        W_18_14         : out    vl_logic;
        W_18_15         : out    vl_logic;
        W_18_16         : out    vl_logic;
        W_18_17         : out    vl_logic;
        W_18_18         : out    vl_logic;
        W_18_19         : out    vl_logic;
        W_18_20         : out    vl_logic;
        W_18_21         : out    vl_logic;
        W_18_22         : out    vl_logic;
        W_18_23         : out    vl_logic;
        W_18_24         : out    vl_logic;
        W_18_25         : out    vl_logic;
        W_18_26         : out    vl_logic;
        W_18_27         : out    vl_logic;
        W_18_28         : out    vl_logic;
        W_18_29         : out    vl_logic;
        W_18_30         : out    vl_logic;
        W_18_31         : out    vl_logic;
        W_17_0          : out    vl_logic;
        W_17_1          : out    vl_logic;
        W_17_2          : out    vl_logic;
        W_17_3          : out    vl_logic;
        W_17_4          : out    vl_logic;
        W_17_5          : out    vl_logic;
        W_17_6          : out    vl_logic;
        W_17_7          : out    vl_logic;
        W_17_8          : out    vl_logic;
        W_17_9          : out    vl_logic;
        W_17_10         : out    vl_logic;
        W_17_11         : out    vl_logic;
        W_17_12         : out    vl_logic;
        W_17_13         : out    vl_logic;
        W_17_14         : out    vl_logic;
        W_17_15         : out    vl_logic;
        W_17_16         : out    vl_logic;
        W_17_17         : out    vl_logic;
        W_17_18         : out    vl_logic;
        W_17_19         : out    vl_logic;
        W_17_20         : out    vl_logic;
        W_17_21         : out    vl_logic;
        W_17_22         : out    vl_logic;
        W_17_23         : out    vl_logic;
        W_17_24         : out    vl_logic;
        W_17_25         : out    vl_logic;
        W_17_26         : out    vl_logic;
        W_17_27         : out    vl_logic;
        W_17_28         : out    vl_logic;
        W_17_29         : out    vl_logic;
        W_17_30         : out    vl_logic;
        W_17_31         : out    vl_logic;
        W_16_0          : out    vl_logic;
        W_16_1          : out    vl_logic;
        W_16_2          : out    vl_logic;
        W_16_3          : out    vl_logic;
        W_16_4          : out    vl_logic;
        W_16_5          : out    vl_logic;
        W_16_6          : out    vl_logic;
        W_16_7          : out    vl_logic;
        W_16_8          : out    vl_logic;
        W_16_9          : out    vl_logic;
        W_16_10         : out    vl_logic;
        W_16_11         : out    vl_logic;
        W_16_12         : out    vl_logic;
        W_16_13         : out    vl_logic;
        W_16_14         : out    vl_logic;
        W_16_15         : out    vl_logic;
        W_16_16         : out    vl_logic;
        W_16_17         : out    vl_logic;
        W_16_18         : out    vl_logic;
        W_16_19         : out    vl_logic;
        W_16_20         : out    vl_logic;
        W_16_21         : out    vl_logic;
        W_16_22         : out    vl_logic;
        W_16_23         : out    vl_logic;
        W_16_24         : out    vl_logic;
        W_16_25         : out    vl_logic;
        W_16_26         : out    vl_logic;
        W_16_27         : out    vl_logic;
        W_16_28         : out    vl_logic;
        W_16_29         : out    vl_logic;
        W_16_30         : out    vl_logic;
        W_16_31         : out    vl_logic;
        W_15_0          : out    vl_logic;
        W_15_1          : out    vl_logic;
        W_15_2          : out    vl_logic;
        W_15_3          : out    vl_logic;
        W_15_4          : out    vl_logic;
        W_15_5          : out    vl_logic;
        W_15_6          : out    vl_logic;
        W_15_7          : out    vl_logic;
        W_15_8          : out    vl_logic;
        W_15_9          : out    vl_logic;
        W_15_10         : out    vl_logic;
        W_15_11         : out    vl_logic;
        W_15_12         : out    vl_logic;
        W_15_13         : out    vl_logic;
        W_15_14         : out    vl_logic;
        W_15_15         : out    vl_logic;
        W_15_16         : out    vl_logic;
        W_15_17         : out    vl_logic;
        W_15_18         : out    vl_logic;
        W_15_19         : out    vl_logic;
        W_15_20         : out    vl_logic;
        W_15_21         : out    vl_logic;
        W_15_22         : out    vl_logic;
        W_15_23         : out    vl_logic;
        W_15_24         : out    vl_logic;
        W_15_25         : out    vl_logic;
        W_15_26         : out    vl_logic;
        W_15_27         : out    vl_logic;
        W_15_28         : out    vl_logic;
        W_15_29         : out    vl_logic;
        W_15_30         : out    vl_logic;
        W_15_31         : out    vl_logic;
        W_14_0          : out    vl_logic;
        W_14_1          : out    vl_logic;
        W_14_2          : out    vl_logic;
        W_14_3          : out    vl_logic;
        W_14_4          : out    vl_logic;
        W_14_5          : out    vl_logic;
        W_14_6          : out    vl_logic;
        W_14_7          : out    vl_logic;
        W_14_8          : out    vl_logic;
        W_14_9          : out    vl_logic;
        W_14_10         : out    vl_logic;
        W_14_11         : out    vl_logic;
        W_14_12         : out    vl_logic;
        W_14_13         : out    vl_logic;
        W_14_14         : out    vl_logic;
        W_14_15         : out    vl_logic;
        W_14_16         : out    vl_logic;
        W_14_17         : out    vl_logic;
        W_14_18         : out    vl_logic;
        W_14_19         : out    vl_logic;
        W_14_20         : out    vl_logic;
        W_14_21         : out    vl_logic;
        W_14_22         : out    vl_logic;
        W_14_23         : out    vl_logic;
        W_14_24         : out    vl_logic;
        W_14_25         : out    vl_logic;
        W_14_26         : out    vl_logic;
        W_14_27         : out    vl_logic;
        W_14_28         : out    vl_logic;
        W_14_29         : out    vl_logic;
        W_14_30         : out    vl_logic;
        W_14_31         : out    vl_logic;
        W_13_0          : out    vl_logic;
        W_13_1          : out    vl_logic;
        W_13_2          : out    vl_logic;
        W_13_3          : out    vl_logic;
        W_13_4          : out    vl_logic;
        W_13_5          : out    vl_logic;
        W_13_6          : out    vl_logic;
        W_13_7          : out    vl_logic;
        W_13_8          : out    vl_logic;
        W_13_9          : out    vl_logic;
        W_13_10         : out    vl_logic;
        W_13_11         : out    vl_logic;
        W_13_12         : out    vl_logic;
        W_13_13         : out    vl_logic;
        W_13_14         : out    vl_logic;
        W_13_15         : out    vl_logic;
        W_13_16         : out    vl_logic;
        W_13_17         : out    vl_logic;
        W_13_18         : out    vl_logic;
        W_13_19         : out    vl_logic;
        W_13_20         : out    vl_logic;
        W_13_21         : out    vl_logic;
        W_13_22         : out    vl_logic;
        W_13_23         : out    vl_logic;
        W_13_24         : out    vl_logic;
        W_13_25         : out    vl_logic;
        W_13_26         : out    vl_logic;
        W_13_27         : out    vl_logic;
        W_13_28         : out    vl_logic;
        W_13_29         : out    vl_logic;
        W_13_30         : out    vl_logic;
        W_13_31         : out    vl_logic;
        W_12_0          : out    vl_logic;
        W_12_1          : out    vl_logic;
        W_12_2          : out    vl_logic;
        W_12_3          : out    vl_logic;
        W_12_4          : out    vl_logic;
        W_12_5          : out    vl_logic;
        W_12_6          : out    vl_logic;
        W_12_7          : out    vl_logic;
        W_12_8          : out    vl_logic;
        W_12_9          : out    vl_logic;
        W_12_10         : out    vl_logic;
        W_12_11         : out    vl_logic;
        W_12_12         : out    vl_logic;
        W_12_13         : out    vl_logic;
        W_12_14         : out    vl_logic;
        W_12_15         : out    vl_logic;
        W_12_16         : out    vl_logic;
        W_12_17         : out    vl_logic;
        W_12_18         : out    vl_logic;
        W_12_19         : out    vl_logic;
        W_12_20         : out    vl_logic;
        W_12_21         : out    vl_logic;
        W_12_22         : out    vl_logic;
        W_12_23         : out    vl_logic;
        W_12_24         : out    vl_logic;
        W_12_25         : out    vl_logic;
        W_12_26         : out    vl_logic;
        W_12_27         : out    vl_logic;
        W_12_28         : out    vl_logic;
        W_12_29         : out    vl_logic;
        W_12_30         : out    vl_logic;
        W_12_31         : out    vl_logic;
        W_11_0          : out    vl_logic;
        W_11_1          : out    vl_logic;
        W_11_2          : out    vl_logic;
        W_11_3          : out    vl_logic;
        W_11_4          : out    vl_logic;
        W_11_5          : out    vl_logic;
        W_11_6          : out    vl_logic;
        W_11_7          : out    vl_logic;
        W_11_8          : out    vl_logic;
        W_11_9          : out    vl_logic;
        W_11_10         : out    vl_logic;
        W_11_11         : out    vl_logic;
        W_11_12         : out    vl_logic;
        W_11_13         : out    vl_logic;
        W_11_14         : out    vl_logic;
        W_11_15         : out    vl_logic;
        W_11_16         : out    vl_logic;
        W_11_17         : out    vl_logic;
        W_11_18         : out    vl_logic;
        W_11_19         : out    vl_logic;
        W_11_20         : out    vl_logic;
        W_11_21         : out    vl_logic;
        W_11_22         : out    vl_logic;
        W_11_23         : out    vl_logic;
        W_11_24         : out    vl_logic;
        W_11_25         : out    vl_logic;
        W_11_26         : out    vl_logic;
        W_11_27         : out    vl_logic;
        W_11_28         : out    vl_logic;
        W_11_29         : out    vl_logic;
        W_11_30         : out    vl_logic;
        W_11_31         : out    vl_logic;
        W_10_0          : out    vl_logic;
        W_10_1          : out    vl_logic;
        W_10_2          : out    vl_logic;
        W_10_3          : out    vl_logic;
        W_10_4          : out    vl_logic;
        W_10_5          : out    vl_logic;
        W_10_6          : out    vl_logic;
        W_10_7          : out    vl_logic;
        W_10_8          : out    vl_logic;
        W_10_9          : out    vl_logic;
        W_10_10         : out    vl_logic;
        W_10_11         : out    vl_logic;
        W_10_12         : out    vl_logic;
        W_10_13         : out    vl_logic;
        W_10_14         : out    vl_logic;
        W_10_15         : out    vl_logic;
        W_10_16         : out    vl_logic;
        W_10_17         : out    vl_logic;
        W_10_18         : out    vl_logic;
        W_10_19         : out    vl_logic;
        W_10_20         : out    vl_logic;
        W_10_21         : out    vl_logic;
        W_10_22         : out    vl_logic;
        W_10_23         : out    vl_logic;
        W_10_24         : out    vl_logic;
        W_10_25         : out    vl_logic;
        W_10_26         : out    vl_logic;
        W_10_27         : out    vl_logic;
        W_10_28         : out    vl_logic;
        W_10_29         : out    vl_logic;
        W_10_30         : out    vl_logic;
        W_10_31         : out    vl_logic;
        W_9_0           : out    vl_logic;
        W_9_1           : out    vl_logic;
        W_9_2           : out    vl_logic;
        W_9_3           : out    vl_logic;
        W_9_4           : out    vl_logic;
        W_9_5           : out    vl_logic;
        W_9_6           : out    vl_logic;
        W_9_7           : out    vl_logic;
        W_9_8           : out    vl_logic;
        W_9_9           : out    vl_logic;
        W_9_10          : out    vl_logic;
        W_9_11          : out    vl_logic;
        W_9_12          : out    vl_logic;
        W_9_13          : out    vl_logic;
        W_9_14          : out    vl_logic;
        W_9_15          : out    vl_logic;
        W_9_16          : out    vl_logic;
        W_9_17          : out    vl_logic;
        W_9_18          : out    vl_logic;
        W_9_19          : out    vl_logic;
        W_9_20          : out    vl_logic;
        W_9_21          : out    vl_logic;
        W_9_22          : out    vl_logic;
        W_9_23          : out    vl_logic;
        W_9_24          : out    vl_logic;
        W_9_25          : out    vl_logic;
        W_9_26          : out    vl_logic;
        W_9_27          : out    vl_logic;
        W_9_28          : out    vl_logic;
        W_9_29          : out    vl_logic;
        W_9_30          : out    vl_logic;
        W_9_31          : out    vl_logic;
        W_8_0           : out    vl_logic;
        W_8_1           : out    vl_logic;
        W_8_2           : out    vl_logic;
        W_8_3           : out    vl_logic;
        W_8_4           : out    vl_logic;
        W_8_5           : out    vl_logic;
        W_8_6           : out    vl_logic;
        W_8_7           : out    vl_logic;
        W_8_8           : out    vl_logic;
        W_8_9           : out    vl_logic;
        W_8_10          : out    vl_logic;
        W_8_11          : out    vl_logic;
        W_8_12          : out    vl_logic;
        W_8_13          : out    vl_logic;
        W_8_14          : out    vl_logic;
        W_8_15          : out    vl_logic;
        W_8_16          : out    vl_logic;
        W_8_17          : out    vl_logic;
        W_8_18          : out    vl_logic;
        W_8_19          : out    vl_logic;
        W_8_20          : out    vl_logic;
        W_8_21          : out    vl_logic;
        W_8_22          : out    vl_logic;
        W_8_23          : out    vl_logic;
        W_8_24          : out    vl_logic;
        W_8_25          : out    vl_logic;
        W_8_26          : out    vl_logic;
        W_8_27          : out    vl_logic;
        W_8_28          : out    vl_logic;
        W_8_29          : out    vl_logic;
        W_8_30          : out    vl_logic;
        W_8_31          : out    vl_logic;
        W_7_0           : out    vl_logic;
        W_7_1           : out    vl_logic;
        W_7_2           : out    vl_logic;
        W_7_3           : out    vl_logic;
        W_7_4           : out    vl_logic;
        W_7_5           : out    vl_logic;
        W_7_6           : out    vl_logic;
        W_7_7           : out    vl_logic;
        W_7_8           : out    vl_logic;
        W_7_9           : out    vl_logic;
        W_7_10          : out    vl_logic;
        W_7_11          : out    vl_logic;
        W_7_12          : out    vl_logic;
        W_7_13          : out    vl_logic;
        W_7_14          : out    vl_logic;
        W_7_15          : out    vl_logic;
        W_7_16          : out    vl_logic;
        W_7_17          : out    vl_logic;
        W_7_18          : out    vl_logic;
        W_7_19          : out    vl_logic;
        W_7_20          : out    vl_logic;
        W_7_21          : out    vl_logic;
        W_7_22          : out    vl_logic;
        W_7_23          : out    vl_logic;
        W_7_24          : out    vl_logic;
        W_7_25          : out    vl_logic;
        W_7_26          : out    vl_logic;
        W_7_27          : out    vl_logic;
        W_7_28          : out    vl_logic;
        W_7_29          : out    vl_logic;
        W_7_30          : out    vl_logic;
        W_7_31          : out    vl_logic;
        W_6_0           : out    vl_logic;
        W_6_1           : out    vl_logic;
        W_6_2           : out    vl_logic;
        W_6_3           : out    vl_logic;
        W_6_4           : out    vl_logic;
        W_6_5           : out    vl_logic;
        W_6_6           : out    vl_logic;
        W_6_7           : out    vl_logic;
        W_6_8           : out    vl_logic;
        W_6_9           : out    vl_logic;
        W_6_10          : out    vl_logic;
        W_6_11          : out    vl_logic;
        W_6_12          : out    vl_logic;
        W_6_13          : out    vl_logic;
        W_6_14          : out    vl_logic;
        W_6_15          : out    vl_logic;
        W_6_16          : out    vl_logic;
        W_6_17          : out    vl_logic;
        W_6_18          : out    vl_logic;
        W_6_19          : out    vl_logic;
        W_6_20          : out    vl_logic;
        W_6_21          : out    vl_logic;
        W_6_22          : out    vl_logic;
        W_6_23          : out    vl_logic;
        W_6_24          : out    vl_logic;
        W_6_25          : out    vl_logic;
        W_6_26          : out    vl_logic;
        W_6_27          : out    vl_logic;
        W_6_28          : out    vl_logic;
        W_6_29          : out    vl_logic;
        W_6_30          : out    vl_logic;
        W_6_31          : out    vl_logic;
        W_5_0           : out    vl_logic;
        W_5_1           : out    vl_logic;
        W_5_2           : out    vl_logic;
        W_5_3           : out    vl_logic;
        W_5_4           : out    vl_logic;
        W_5_5           : out    vl_logic;
        W_5_6           : out    vl_logic;
        W_5_7           : out    vl_logic;
        W_5_8           : out    vl_logic;
        W_5_9           : out    vl_logic;
        W_5_10          : out    vl_logic;
        W_5_11          : out    vl_logic;
        W_5_12          : out    vl_logic;
        W_5_13          : out    vl_logic;
        W_5_14          : out    vl_logic;
        W_5_15          : out    vl_logic;
        W_5_16          : out    vl_logic;
        W_5_17          : out    vl_logic;
        W_5_18          : out    vl_logic;
        W_5_19          : out    vl_logic;
        W_5_20          : out    vl_logic;
        W_5_21          : out    vl_logic;
        W_5_22          : out    vl_logic;
        W_5_23          : out    vl_logic;
        W_5_24          : out    vl_logic;
        W_5_25          : out    vl_logic;
        W_5_26          : out    vl_logic;
        W_5_27          : out    vl_logic;
        W_5_28          : out    vl_logic;
        W_5_29          : out    vl_logic;
        W_5_30          : out    vl_logic;
        W_5_31          : out    vl_logic;
        W_4_0           : out    vl_logic;
        W_4_1           : out    vl_logic;
        W_4_2           : out    vl_logic;
        W_4_3           : out    vl_logic;
        W_4_4           : out    vl_logic;
        W_4_5           : out    vl_logic;
        W_4_6           : out    vl_logic;
        W_4_7           : out    vl_logic;
        W_4_8           : out    vl_logic;
        W_4_9           : out    vl_logic;
        W_4_10          : out    vl_logic;
        W_4_11          : out    vl_logic;
        W_4_12          : out    vl_logic;
        W_4_13          : out    vl_logic;
        W_4_14          : out    vl_logic;
        W_4_15          : out    vl_logic;
        W_4_16          : out    vl_logic;
        W_4_17          : out    vl_logic;
        W_4_18          : out    vl_logic;
        W_4_19          : out    vl_logic;
        W_4_20          : out    vl_logic;
        W_4_21          : out    vl_logic;
        W_4_22          : out    vl_logic;
        W_4_23          : out    vl_logic;
        W_4_24          : out    vl_logic;
        W_4_25          : out    vl_logic;
        W_4_26          : out    vl_logic;
        W_4_27          : out    vl_logic;
        W_4_28          : out    vl_logic;
        W_4_29          : out    vl_logic;
        W_4_30          : out    vl_logic;
        W_4_31          : out    vl_logic;
        W_3_0           : out    vl_logic;
        W_3_1           : out    vl_logic;
        W_3_2           : out    vl_logic;
        W_3_3           : out    vl_logic;
        W_3_4           : out    vl_logic;
        W_3_5           : out    vl_logic;
        W_3_6           : out    vl_logic;
        W_3_7           : out    vl_logic;
        W_3_8           : out    vl_logic;
        W_3_9           : out    vl_logic;
        W_3_10          : out    vl_logic;
        W_3_11          : out    vl_logic;
        W_3_12          : out    vl_logic;
        W_3_13          : out    vl_logic;
        W_3_14          : out    vl_logic;
        W_3_15          : out    vl_logic;
        W_3_16          : out    vl_logic;
        W_3_17          : out    vl_logic;
        W_3_18          : out    vl_logic;
        W_3_19          : out    vl_logic;
        W_3_20          : out    vl_logic;
        W_3_21          : out    vl_logic;
        W_3_22          : out    vl_logic;
        W_3_23          : out    vl_logic;
        W_3_24          : out    vl_logic;
        W_3_25          : out    vl_logic;
        W_3_26          : out    vl_logic;
        W_3_27          : out    vl_logic;
        W_3_28          : out    vl_logic;
        W_3_29          : out    vl_logic;
        W_3_30          : out    vl_logic;
        W_3_31          : out    vl_logic;
        W_2_0           : out    vl_logic;
        W_2_1           : out    vl_logic;
        W_2_2           : out    vl_logic;
        W_2_3           : out    vl_logic;
        W_2_4           : out    vl_logic;
        W_2_5           : out    vl_logic;
        W_2_6           : out    vl_logic;
        W_2_7           : out    vl_logic;
        W_2_8           : out    vl_logic;
        W_2_9           : out    vl_logic;
        W_2_10          : out    vl_logic;
        W_2_11          : out    vl_logic;
        W_2_12          : out    vl_logic;
        W_2_13          : out    vl_logic;
        W_2_14          : out    vl_logic;
        W_2_15          : out    vl_logic;
        W_2_16          : out    vl_logic;
        W_2_17          : out    vl_logic;
        W_2_18          : out    vl_logic;
        W_2_19          : out    vl_logic;
        W_2_20          : out    vl_logic;
        W_2_21          : out    vl_logic;
        W_2_22          : out    vl_logic;
        W_2_23          : out    vl_logic;
        W_2_24          : out    vl_logic;
        W_2_25          : out    vl_logic;
        W_2_26          : out    vl_logic;
        W_2_27          : out    vl_logic;
        W_2_28          : out    vl_logic;
        W_2_29          : out    vl_logic;
        W_2_30          : out    vl_logic;
        W_2_31          : out    vl_logic;
        W_1_0           : out    vl_logic;
        W_1_1           : out    vl_logic;
        W_1_2           : out    vl_logic;
        W_1_3           : out    vl_logic;
        W_1_4           : out    vl_logic;
        W_1_5           : out    vl_logic;
        W_1_6           : out    vl_logic;
        W_1_7           : out    vl_logic;
        W_1_8           : out    vl_logic;
        W_1_9           : out    vl_logic;
        W_1_10          : out    vl_logic;
        W_1_11          : out    vl_logic;
        W_1_12          : out    vl_logic;
        W_1_13          : out    vl_logic;
        W_1_14          : out    vl_logic;
        W_1_15          : out    vl_logic;
        W_1_16          : out    vl_logic;
        W_1_17          : out    vl_logic;
        W_1_18          : out    vl_logic;
        W_1_19          : out    vl_logic;
        W_1_20          : out    vl_logic;
        W_1_21          : out    vl_logic;
        W_1_22          : out    vl_logic;
        W_1_23          : out    vl_logic;
        W_1_24          : out    vl_logic;
        W_1_25          : out    vl_logic;
        W_1_26          : out    vl_logic;
        W_1_27          : out    vl_logic;
        W_1_28          : out    vl_logic;
        W_1_29          : out    vl_logic;
        W_1_30          : out    vl_logic;
        W_1_31          : out    vl_logic;
        W_0_0           : out    vl_logic;
        W_0_1           : out    vl_logic;
        W_0_2           : out    vl_logic;
        W_0_3           : out    vl_logic;
        W_0_4           : out    vl_logic;
        W_0_5           : out    vl_logic;
        W_0_6           : out    vl_logic;
        W_0_7           : out    vl_logic;
        W_0_8           : out    vl_logic;
        W_0_9           : out    vl_logic;
        W_0_10          : out    vl_logic;
        W_0_11          : out    vl_logic;
        W_0_12          : out    vl_logic;
        W_0_13          : out    vl_logic;
        W_0_14          : out    vl_logic;
        W_0_15          : out    vl_logic;
        W_0_16          : out    vl_logic;
        W_0_17          : out    vl_logic;
        W_0_18          : out    vl_logic;
        W_0_19          : out    vl_logic;
        W_0_20          : out    vl_logic;
        W_0_21          : out    vl_logic;
        W_0_22          : out    vl_logic;
        W_0_23          : out    vl_logic;
        W_0_24          : out    vl_logic;
        W_0_25          : out    vl_logic;
        W_0_26          : out    vl_logic;
        W_0_27          : out    vl_logic;
        W_0_28          : out    vl_logic;
        W_0_29          : out    vl_logic;
        W_0_30          : out    vl_logic;
        W_0_31          : out    vl_logic
    );
end MessageScheduler;
